module alutest(input[15:0] a,b,input[3:0] switch,output[15:0] op);
	wire [15:0]sumxy,diffxy,diffyx,r0,r1,rn1,negx,negy,xbar,ybar,xin,yin,xde,yde,xandy,xory;
    addsub a1(sumxy,a,b,1'b0);
   	addsub a2(diffxy,a,b,1'b1);
  	addsub a3(diffyx,b,a,1'b1);
  	addsub z1(r0,16'b0,16'b0,1'b0);
  	addsub o1(r1,16'b0,0000000000000001,1'b0);
  	addsub m1(rn1,16'b0,0000000000000001,1'b1);
  	addsub a4(negx,16'b0,a,1'b1);
  	addsub a5(negy,16'b0,b,1'b1);
	negator n1(xbar,a);
	negator n2(ybar,b);
  	addsub a6(xin,a,0000000000000001,1'b0);
  	addsub a7(yin,b,0000000000000001,1'b0);
  	addsub s8(xde,a,0000000000000001,1'b1);
  	addsub s9(yde,b,0000000000000001,1'b1);
	andop aop1(xandy,a,b);
	orop oop1(xory,a,b);
	mux m2(op,switch,sumxy,diffxy,diffyx,r0,r1,rn1,negx,negy,xbar,ybar,xin,yin,xde,yde,xandy,xory);
endmodule
module andop(output[15:0] c,input[15:0]a,b);
	and_gate a0(c[0],a[0],b[0]);
	and_gate a1(c[1],a[1],b[1]);
	and_gate a2(c[2],a[2],b[2]);
	and_gate a3(c[3],a[3],b[3]);
	and_gate a4(c[4],a[4],b[4]);
	and_gate a5(c[5],a[5],b[5]);
	and_gate a6(c[6],a[6],b[6]);
	and_gate a7(c[7],a[7],b[7]);
	and_gate a8(c[8],a[8],b[8]);
	and_gate a9(c[9],a[9],b[9]);
	and_gate a10(c[10],a[10],b[10]);
	and_gate a11(c[11],a[11],b[11]);
	and_gate a12(c[12],a[12],b[12]);
	and_gate a13(c[13],a[13],b[13]);
	and_gate a14(c[14],a[14],b[14]);
	and_gate a15(c[15],a[15],b[15]);
endmodule
module orop(output[15:0] c,input[15:0]a,b);
	or_gate a0(c[0],a[0],b[0]);
	or_gate a1(c[1],a[1],b[1]);
	or_gate a2(c[2],a[2],b[2]);
	or_gate a3(c[3],a[3],b[3]);
	or_gate a4(c[4],a[4],b[4]);
	or_gate a5(c[5],a[5],b[5]);
	or_gate a6(c[6],a[6],b[6]);
	or_gate a7(c[7],a[7],b[7]);
	or_gate a8(c[8],a[8],b[8]);
	or_gate a9(c[9],a[9],b[9]);
	or_gate a10(c[10],a[10],b[10]);
	or_gate a11(c[11],a[11],b[11]);
	or_gate a12(c[12],a[12],b[12]);
	or_gate a13(c[13],a[13],b[13]);
	or_gate a14(c[14],a[14],b[14]);
	or_gate a15(c[15],a[15],b[15]);
endmodule
module negator(output[15:0] b,input[15:0] a);
	notgate n0(b[0],a[0]);
	notgate n1(b[1],a[1]);
	notgate n2(b[2],a[2]);
	notgate n3(b[3],a[3]);
	notgate n4(b[4],a[4]);
	notgate n5(b[5],a[5]);
	notgate n6(b[6],a[6]);
	notgate n7(b[7],a[7]);
	notgate n8(b[8],a[8]);
	notgate n9(b[9],a[9]);
	notgate n10(b[10],a[10]);	
	notgate n11(b[11],a[11]);
	notgate n12(b[12],a[12]);
	notgate n13(b[13],a[13]);
	notgate n14(b[14],a[14]);
	notgate n15(b[15],a[15]);
endmodule
module addsub(s,a,b,m);
  	input [15:0]a,b;
  	input m;
	output [15:0]s;
  	wire [15:0]c;
  	wire [15:0] var1;
  	xor_gate x0(var1[0],b[0],m);
  	xor_gate x1(var1[1],b[1],m);
  	xor_gate x2(var1[2],b[2],m);
  	xor_gate x3(var1[3],b[3],m);
  	xor_gate x4(var1[4],b[4],m);
  	xor_gate x5(var1[5],b[5],m);
  	xor_gate x6(var1[6],b[6],m);
  	xor_gate x7(var1[7],b[7],m);
  	xor_gate x8(var1[8],b[8],m);
  	xor_gate x9(var1[9],b[9],m);
  	xor_gate x10(var1[10],b[10],m);
  	xor_gate x11(var1[11],b[11],m);
  	xor_gate x12(var1[12],b[12],m);
  	xor_gate x13(var1[13],b[13],m);
  	xor_gate x14(var1[14],b[14],m);
  	xor_gate x15(var1[15],b[15],m);
  	full f0(s[0],c[0],a[0],var1[0],m);
  	full f1(s[1],c[1],a[1],var1[1],c[0]);
  	full f2(s[2],c[2],a[2],var1[2],c[1]);
  	full f3(s[3],c[3],a[3],var1[3],c[2]);
  	full f4(s[4],c[4],a[4],var1[4],c[3]);
  	full f5(s[5],c[5],a[5],var1[5],c[4]);
  	full f6(s[6],c[6],a[6],var1[6],c[5]);
  	full f7(s[7],c[7],a[7],var1[7],c[6]);
  	full f8(s[8],c[8],a[8],var1[8],c[7]);
  	full f9(s[9],c[9],a[9],var1[9],c[8]);
  	full f10(s[10],c[10],a[10],var1[10],c[9]);
  	full f11(s[11],c[11],a[11],var1[11],c[10]);
  	full f12(s[12],c[12],a[12],var1[12],c[11]);
  	full f13(s[13],c[13],a[13],var1[13],c[12]);
  	full f14(s[14],c[14],a[14],var1[14],c[13]);
  	full f15(s[15],c[15],a[15],var1[15],c[14]);
endmodule
module full(s,c,a,b,d);
  	input a,b,d;
  	output s,c;
  	wire s1,c1,c2;
  	half h0(s1,c1,a,b);
  	half h1(s,c2,s1,d);
  	or_gate o1(c,c1,c2);
endmodule
module half(s,c,a,b);
  	input a,b;
  	output s,c;
  	xor_gate x1(s,a,b);
  	and_gate a1(c,a,b);
endmodule
module or_gate(output c,input a,b);
	wire x;
	nor(x,a,b);
	nor(c,x,x);
endmodule
module notgate(output b,input a);
	nand(b,a,a);
endmodule
module and_gate(output c,input a,b);
	wire x;
	nand(x,a,b);
	nand(c,x,x);
endmodule
module xor_gate(output c,input a,b);
	wire x,y,z;
	nand(x,a,b);
	nand(y,a,x);
	nand(z,b,x);
	nand(c,y,z);
endmodule
module mux(output[15:0]op,input[3:0] s,input[16:0]a,b,c,d,e,f,g,h,i,j,k,l,m,n,o,p);
	wire[3:0] sn;
	wire[16:0] at,bt,ct,dt,et,ft,gt,ht,it,jt,kt,lt,mt,nt,ot,pt;
	wire[16:0]check;
  	notgate n0(sn[0],s[0]);
  	notgate n1(sn[1],s[1]);
	notgate n2(sn[2],s[2]);
	notgate n3(sn[3],s[3]);
  	submux s0(at,a,sn[3],sn[2],sn[1],sn[0]);
  	submux s1(bt,b,sn[3],sn[2],sn[1],s[0]);
  	submux s2(ct,c,sn[3],sn[2],s[1],sn[0]);
  	submux s3(dt,d,sn[3],sn[2],s[1],s[0]);
  	submux s4(et,e,sn[3],s[2],sn[1],sn[0]);
  	submux s5(ft,f,sn[3],s[2],sn[1],s[0]);
  	submux s6(gt,g,sn[3],s[2],s[1],sn[0]);
  	submux s7(ht,h,sn[3],s[2],s[1],s[0]);
  	submux s8(it,i,s[3],sn[2],sn[1],sn[0]);
  	submux s9(jt,j,s[3],sn[2],sn[1],s[0]);
  	submux s10(kt,k,s[3],sn[2],s[1],sn[0]);
  	submux s11(lt,l,s[3],sn[2],s[1],s[0]);
  	submux s12(mt,m,s[3],s[2],sn[1],sn[0]);
  	submux s13(nt,n,s[3],s[2],sn[1],s[0]);
  	submux s14(ot,o,s[3],s[2],s[1],sn[0]);
  	submux s15(pt,p,s[3],s[2],s[1],s[0]);
	or16bit o0(op[0],at[0],bt[0],ct[0],dt[0],et[0],ft[0],gt[0],ht[0],it[0],jt[0],kt[0],lt[0],mt[0],nt[0],ot[0],pt[0]);
	or16bit o1(op[1],at[1],bt[1],ct[1],dt[1],et[1],ft[1],gt[1],ht[1],it[1],jt[1],kt[1],lt[1],mt[1],nt[1],ot[1],pt[1]);
	or16bit o2(op[2],at[2],bt[2],ct[2],dt[2],et[2],ft[2],gt[2],ht[2],it[2],jt[2],kt[2],lt[2],mt[2],nt[2],ot[2],pt[2]);
	or16bit o3(op[3],at[3],bt[3],ct[3],dt[3],et[3],ft[3],gt[3],ht[3],it[3],jt[3],kt[3],lt[3],mt[3],nt[3],ot[3],pt[3]);
	or16bit o4(op[4],at[4],bt[4],ct[4],dt[4],et[4],ft[4],gt[4],ht[4],it[4],jt[4],kt[4],lt[4],mt[4],nt[4],ot[4],pt[4]);
	or16bit o5(op[5],at[5],bt[5],ct[5],dt[5],et[5],ft[5],gt[5],ht[5],it[5],jt[5],kt[5],lt[5],mt[5],nt[5],ot[5],pt[5]);
	or16bit o6(op[6],at[6],bt[6],ct[6],dt[6],et[6],ft[6],gt[6],ht[6],it[6],jt[6],kt[6],lt[6],mt[6],nt[6],ot[6],pt[6]);
	or16bit o7(op[7],at[7],bt[7],ct[7],dt[7],et[7],ft[7],gt[7],ht[7],it[7],jt[7],kt[7],lt[7],mt[7],nt[7],ot[7],pt[7]);
	or16bit o8(op[8],at[8],bt[8],ct[8],dt[8],et[8],ft[8],gt[8],ht[8],it[8],jt[8],kt[8],lt[8],mt[8],nt[8],ot[8],pt[8]);
	or16bit o9(op[9],at[9],bt[9],ct[9],dt[9],et[9],ft[9],gt[9],ht[9],it[9],jt[9],kt[9],lt[9],mt[9],nt[9],ot[9],pt[9]);
	or16bit o10(op[10],at[10],bt[10],ct[10],dt[10],et[10],ft[10],gt[10],ht[10],it[10],jt[10],kt[10],lt[10],mt[10],nt[10],ot[10],pt[10]);
	or16bit o11(op[11],at[11],bt[11],ct[11],dt[11],et[11],ft[11],gt[11],ht[11],it[11],jt[11],kt[11],lt[11],mt[11],nt[11],ot[11],pt[11]);
	or16bit o12(op[12],at[12],bt[12],ct[12],dt[12],et[12],ft[12],gt[12],ht[12],it[12],jt[12],kt[12],lt[12],mt[12],nt[12],ot[12],pt[12]);
	or16bit o13(op[13],at[13],bt[13],ct[13],dt[13],et[13],ft[13],gt[13],ht[13],it[13],jt[13],kt[13],lt[13],mt[13],nt[13],ot[13],pt[13]);
	or16bit o14(op[14],at[14],bt[14],ct[14],dt[14],et[14],ft[14],gt[14],ht[14],it[14],jt[14],kt[14],lt[14],mt[14],nt[14],ot[14],pt[14]);
	or16bit o15(op[15],at[15],bt[15],ct[15],dt[15],et[15],ft[15],gt[15],ht[15],it[15],jt[15],kt[15],lt[15],mt[15],nt[15],ot[15],pt[15]);
endmodule
module submux(output[15:0] op,input[15:0] a,input b,c,d,e);
	and5gate a0(op[0],a[0],b,c,d,e);
	and5gate a1(op[1],a[1],b,c,d,e);
	and5gate a2(op[2],a[2],b,c,d,e);
	and5gate a3(op[3],a[3],b,c,d,e);
	and5gate a4(op[4],a[4],b,c,d,e);
	and5gate a5(op[5],a[5],b,c,d,e);
	and5gate a6(op[6],a[6],b,c,d,e);
	and5gate a7(op[7],a[7],b,c,d,e);
	and5gate a8(op[8],a[8],b,c,d,e);
	and5gate a9(op[9],a[9],b,c,d,e);
	and5gate a10(op[10],a[10],b,c,d,e);
	and5gate a11(op[11],a[11],b,c,d,e);
	and5gate a12(op[12],a[12],b,c,d,e);
	and5gate a13(op[13],a[13],b,c,d,e);
	and5gate a14(op[14],a[14],b,c,d,e);
	and5gate a15(op[15],a[15],b,c,d,e);
endmodule
module and5gate(output op,input a,b,c,d,e);
	wire p,q,r;
	and_gate a0(p,a,b);
	and_gate a1(q,p,c);
	and_gate a2(r,q,d);
	and_gate a3(op,r,e);
endmodule
module or16bit(output op,input i1,i2,i3,i4,i5,i6,i7,i8,j1,j2,j3,j4,j5,j6,j7,j8);
	wire a,b,c,d,e,f,g,h,i,j,k,l,m,n;
	or_gate o0(a,i1,i2);
	or_gate o1(b,a,i3);
	or_gate o2(c,b,i4);
	or_gate o3(d,c,i5);
	or_gate o4(e,d,i6);
	or_gate o5(f,e,i7);
	or_gate o6(g,f,i8);
	or_gate o7(h,g,j1);
	or_gate o8(i,h,j2);
	or_gate o9(j,i,j3);
	or_gate o10(k,j,j4);
	or_gate o11(l,k,j5);
	or_gate o12(m,l,j6);
	or_gate o13(n,m,j7);
	or_gate o14(op,n,j8);
endmodule

module alutest_test;
	reg[15:0] a,b;
	reg[3:0] switch;
	wire[15:0] op;
	alutest test(a,b,switch,op);
	integer count;
	initial begin
  		$dumpfile("dump.vcd");
  		$dumpvars;
  		a={$random}%65536;
  		b={$random}%65536;
		for(count=0;count<16;count=count+1)begin
			{switch}=count;
			#20;
		end
	end
endmodule
